`timescale 1ns / 1ns 
module ha_tb;

reg a, b;
wire sum, cout;
integer i;

ha ha_DUT (.a(a), .b(b), .sum(sum), .cout(cout));

initial begin

#10
a <= 0; b <= 0;

for (i = 0; i < 4; i = i + 1) begin
	
	{a, b} = i;
	#10;
	
end

$stop;

end

endmodule