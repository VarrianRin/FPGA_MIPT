`timescale 1ns / 1ns 
module mux_2x1_tb;

reg a, b, sel;
wire c;
integer i;

mux_2x1 mux_2x1_DUT (.a(a), .b(b), .sel(sel), .c(c));

initial begin

#10
a <= 0; b <= 0; sel <= 0;

for (i = 0; i < 3; i = i + 1) begin
	
	{a, b, sel} = i;
	#10;
	
end

$stop;

end

endmodule