`timescale 1ns / 1ns 
module combo_tb;

reg a, b, c, d;
wire o;

combo combo_DUT (.a(a), .b(b), .c(c), .d(d), .o(o));

initial begin

#10
a = 0; b = 0; c = 0; d = 0;

#10
a = 1; b = 0; c = 0; d = 0;

#10
a = 0; b = 1; c = 0; d = 0;

#10
a = 1; b = 1; c = 0; d = 0;

#10
a = 0; b = 0; c = 1; d = 0;

#10
a = 1; b = 0; c = 1; d = 0;

#10
a = 0; b = 1; c = 1; d = 0;

#10
a = 1; b = 1; c = 1; d = 0;

#10
a = 0; b = 0; c = 0; d = 1;

#10
a = 1; b = 0; c = 0; d = 1;

#10
a = 0; b = 1; c = 0; d = 1;

#10
a = 1; b = 1; c = 0; d = 1;

#10
a = 0; b = 0; c = 1; d = 1;

#10
a = 1; b = 0; c = 1; d = 1;

#10
a = 0; b = 1; c = 1; d = 1;

#10
a = 1; b = 1; c = 1; d = 1;

#10
$stop;

end

endmodule